module Q5_6_1_SDV	(input wire A, B, C, output F);
	
	
endmodule