module Timing(input in, output out);
	assign out = !in;
endmodule