module my_and(input wire A, B, C, output wire F);
	assign F = A & B & C;
endmodule