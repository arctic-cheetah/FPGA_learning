module my_not (input wire A, output wire F);
	assign F = ~A;
endmodule