module first_upload(input in, output out);
	assign out = in;
endmodule